`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:51:17 02/18/2011 
// Design Name: 
// Module Name:    ethernet_clock 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Generate 125 MHz clock 
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ethernet_clock(
    );


endmodule
